`timescale 1ns / 100ps
module mux_tb();
 reg [4:0] ctrl_read;
 reg [31:0] w_0, w_1, w_2, w_3, w_4,
              w_5, w_6, w_7, w_8, w_9, w_10,
				  w_11, w_12, w_13, w_14, w_15,
				  w_16, w_17, w_18, w_19, w_20,
				  w_21, w_22, w_23, w_24, w_25,
				  w_26, w_27, w_28, w_29, w_30, w_31;
 wire [31:0] out;
 
endmodule